module aeqb2 (
    input logic [1:0] a,
    input logic [1:0] b,
    output logic aeqb
);

    /*

     a     b   | aeqb
    -----------+-----
    0 0   0 0  |  1
    0 0   0 1  |  0
    0 0   1 0  |  0
    0 0   1 1  |  0
    0 1   0 0  |  0 
    0 1   0 1  |  1
    0 1   1 0  |  0
    0 1   1 1  |  0
    1 0   0 0  |  0
    1 0   0 1  |  0
    1 0   1 0  |  1
    1 0   1 1  |  0
    1 1   0 0  |  0
    1 1   0 1  |  0
    1 1   1 0  |  0
    1 1   1 1  |  1
    
    */
    
    assign aeqb =
        (~a[1] & ~a[0] & ~b[1] & ~b[0]) |
        (~a[1] &  a[0] & ~b[1] &  b[0]) |
        ( a[1] & ~a[0] &  b[1] & ~b[0]) |
        ( a[1] &  a[0] &  b[1] &  b[0]) ;

endmodule