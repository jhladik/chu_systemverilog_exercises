module agtb2 (
    input logic [1:0] a,
    input logic [1:0] b,
    output logic agtb
);

    /*

     a     b   | agtb
    -----------+-----
    0 0   0 0  |  0
    0 0   0 1  |  0
    0 0   1 0  |  0
    0 0   1 1  |  0
    0 1   0 0  |  1 
    0 1   0 1  |  0
    0 1   1 0  |  0
    0 1   1 1  |  0
    1 0   0 0  |  1
    1 0   0 1  |  1
    1 0   1 0  |  0
    1 0   1 1  |  0
    1 1   0 0  |  1
    1 1   0 1  |  1
    1 1   1 0  |  1
    1 1   1 1  |  0
    
    */
    
    assign agtb =
        (~a[1] &  a[0] & ~b[1] & ~b[0]) |
        ( a[1] & ~a[0] & ~b[1] & ~b[0]) |
        ( a[1] & ~a[0] & ~b[1] &  b[0]) |
        ( a[1] &  a[0] & ~b[1] & ~b[0]) |
        ( a[1] &  a[0] & ~b[1] &  b[0]) |
        ( a[1] &  a[0] &  b[1] & ~b[0]) ;

endmodule